`timescale 1ns / 1ps


module top_uart_fnd(
    input clk,
    input reset,
    input btnr,
    input btnu,
    output [3:0] fndCom,
    output [7:0] fndFont
    );

    
endmodule
